parameter AXI_DATA_WIDTH = 32;
parameter AXI_ADDR_WIDTH = 32;
parameter AXI_STRB_WIDTH = (AXI_DATA_WIDTH+7)/8;

